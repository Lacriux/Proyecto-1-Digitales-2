
module test(
	//--------- Outputs ---------
	output not_a,
	//--------- Inputs ---------
	input a
	
);
	assign not_a = !a;

endmodule
